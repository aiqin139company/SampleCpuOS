module ROM( clk, addr, data );
	input clk;
	input addr;
	output data;
	
	
endmodule
