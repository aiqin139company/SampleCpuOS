module Control_Center( clk, indat, outdat);
	input clk;
	input indat;
	output outdat;
	
endmodule
