module ALU( clk, indat, outdat );
	input clk;
	input indat;
	output outdat;
	
	
endmodule
