module RAM( clk, addr, data);
	input clk;
	input addr;
	inout data;
	
	
endmodule

